�� sr up.mi.jgm.test.CatalogTaǚ#�<b I compteurL relationTabt Ljava/util/ArrayList;xp    sr java.util.ArrayListx����a� I sizexp    w    x