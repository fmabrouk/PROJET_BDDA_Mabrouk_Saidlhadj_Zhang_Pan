�� sr up.mi.jgm.TP04.Catalog\RIo/ � I compteurL Datat Ljava/util/ArrayList;L relationTabq ~ xp    psr java.util.ArrayListx����a� I sizexp   w   sr up.mi.jgm.TP04.RelationInfo��pY19�J L Dataq ~ L nomRelationt Ljava/lang/String;xpsq ~    w   sr up.mi.jgm.TP04.ColInfo�m�A�� I tailleL nomq ~ L typeq ~ xp    t Notest REALsq ~ 	   t Nomt VARCHARxt 	Matièresx